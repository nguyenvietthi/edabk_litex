module neuron_grid_datapath_1x1 #(
    parameter CORE_NUMBER = 0
)(
    input update_potential,
    input local_buffers_full,
    input [255:0] axon_spikes,
    input clk,
    input reset_n,
    input initial_axon_num,
    input inc_axon_num,
    input initial_neuron_num,
    input inc_neuron_num,
    input new_neuron,
    input process_spike,
    output reg done_neuron,
    output done_axon,
    output reg [29:0] packet_out,
    output reg spike_out_valid
);
reg [367:0] neuron_parameter [0:255];
wire [1:0] neuron_instructions[0:255];

wire spike_out;
reg [7:0] axon_num, neuron_num;
wire [8:0] potential_out;


always @(negedge clk, negedge reset_n) begin
    if(~reset_n) begin
        packet_out <= 30'd0;
        spike_out_valid <= 0;
    end
    else begin
        packet_out <= spike_out & update_potential ? neuron_parameter[neuron_num][29:0] : {30{1'b0}};
        spike_out_valid <= (~local_buffers_full) & spike_out & update_potential;
    end
end




assign done_axon = (axon_num == 255);

always @(negedge clk, negedge reset_n) begin
    if(~reset_n) axon_num <= 8'd0;
    else if(initial_axon_num) axon_num <= 8'd0;
    else if(inc_axon_num) axon_num <= axon_num + 1'b1;
    else axon_num <= axon_num;
end

always @(negedge clk, negedge reset_n) begin
    if(~reset_n) neuron_num <= 8'd0;
    else if(initial_neuron_num) neuron_num <= 8'd0;
    else if(inc_neuron_num) neuron_num <= neuron_num + 1'b1;
    else neuron_num <= neuron_num;
end


always @(posedge clk, negedge reset_n) begin
    if(~reset_n) done_neuron <= 0;
    else if(neuron_num == 255) done_neuron <= 1;
    else done_neuron <= 0;
end

wire reg_en;
assign reg_en = (neuron_parameter[neuron_num][112 + axon_num] & axon_spikes[axon_num]);
neuron_block neuron_block(
    .clk(clk),
    .reset_n(reset_n),
    .leak(neuron_parameter[neuron_num][57:49]),
    .weights(neuron_parameter[neuron_num][93:58]),
    .positive_threshold(neuron_parameter[neuron_num][48:40]),
    .negative_threshold(neuron_parameter[neuron_num][39:31]),
    .reset_potential(neuron_parameter[neuron_num][102:94]),
    .current_potential(neuron_parameter[neuron_num][111:103]),
    .neuron_instruction(neuron_instructions[axon_num]),
    .reset_mode(neuron_parameter[neuron_num][30]),
    .new_neuron(new_neuron),
    .process_spike(process_spike),
    .reg_en(reg_en),
    .potential_out(potential_out),
    .spike_out(spike_out)
);

///////Khởi tạo csram
generate
    if(CORE_NUMBER == 0) begin // x = 0, y = 0
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
            neuron_parameter[0] <= 368'b11101010101011111110101010101010001010010010101100000000001010110011010011011010100100100101011101010010101001101101001010010010110110101000011010011110110001111001010001000011100010100010001110111010010100000010101101101010101010101010110001110100011001110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000000000000;
neuron_parameter[1] <= 368'b10011010101110100010101010101001011000001010001110101010101010101101000001011011110100010100101110101001010010111000100100001010100110010000111010100001001011101010100110101111101010101010111010001010101010110001001100001010001000000010100110100101101101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000000010000;
neuron_parameter[2] <= 368'b11101010101011000010010010101001010101011010011101010100000011001101011001011101010100100101100001010000010101101101000000110010010110001001001111011010100101101011101011010111101000110101011010101001010101000010000101010010111010010101001001100101100010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000000100000;
neuron_parameter[3] <= 368'b00001010101011100110111011010010001111011111010110011101011000100001000101101100101001000010110110000110101011011010001100101111101001011010101000101101111010001010101011011011101010101101011010101001010100101011110101010011101010001110111001001110100110010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000000110000;
neuron_parameter[4] <= 368'b00101010101000101110100010101000010000001010101001010000101000100011010010010000100001001001011110100000110010111010011011000111100001101000001110100110101000101011011010000111101101101011001110010010100001100101001100001001001010101010100001100110100101010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000001000000;
neuron_parameter[5] <= 368'b01101010101010010001001001000101110101000000001101010010000000110101000010101100110000101010101010000010101010110001000010101010101000100111011100101010110111100110101011000011111010000100101001010101000110111101010100101001101100001010111110111111111011100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000001010000;
neuron_parameter[6] <= 368'b10101010100011010010101010101001101001001010100110010000010010101001000001001010110000000100101011110110010110110011001001011011101111100100101110101010011010111010101000101011011000001010101010000010101010000001000010100001110101110111011100111010011011000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000001100000;
neuron_parameter[7] <= 368'b01011100010001100010101100100100101010100111011011101010011000110010101000001011101010100100101100100001010000110111000100101011101010001010100000101000101010010010011010011000001101000101000110101100010100000010101010101001011010101010101001110010000010110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000001110000;
neuron_parameter[8] <= 368'b01001010101011001110001000101010101010010010111100101000111011100010000001101011101001000110101110101000001010111010101100101011101010010000111000100100010001101010011011011011001001101000001111001010000110110110100000101011001011101010111111110001110000100000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001000010000000;
neuron_parameter[9] <= 368'b00000101010111011001000101010100100110100101001110001011101110100100101010100010101010110100101010110111010010101011010101101111100101011010011110110100101011101010100010000011101001010100101010100000101010000010101010101011001010101010100100100110111110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000010010000;
neuron_parameter[10] <= 368'b11001010101000110010101010101010001010110100101110100001010010101010100011001011100001101001001010010010100000111001101010000010110000101001001010000010100010101001001000110010000001001000101010100001001010001010110000101010101010101010111010010100010111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000010100000;
neuron_parameter[11] <= 368'b10101010101010110110101010101011011101010000001011110101000101110101010001101011110100100100101110101010000010110000100100101011001011011011011110100101101010111010100010101111101000100111111010101001010100110010000101011010101010100010001101000100111010100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000010110000;
neuron_parameter[12] <= 368'b11101010101011111010010110101011110101001011011011010100101111100101011010001010010100000100101101010001010101111101100010011111010111101011101010110010100101101011011010010110101110110101001010101001010100101010101101010000101010010100001001010111101110100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000011000000;
neuron_parameter[13] <= 368'b11101010101010110110101001010110001010011101010000100010101001000010010010101101101100001010110110111010010010001010100101001011001010101010101010100010101011001011010000010100001000010101011000100000010101110010101010110111101010101010101001010110011001010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000011010000;
neuron_parameter[14] <= 368'b10001010101010101000001001001010001100000100101110000000101010110010100010101111101010010101011110101001000101110010100100010111101000000000101110110000010010101001010000100011100101001010001010010100100000111101001010001011001010101010100011011010111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000011100000;
neuron_parameter[15] <= 368'b11101010101010101110101011001000101010011100111010101101010001110010110000010001101001001010111010111000101010111010101110101110101010100100101111001011010010101101101100001011110000111010101100010010001010110101111001101001101011101010100110001110010111110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000011110000;
neuron_parameter[16] <= 368'b10101010101000100110101010101011101010000010100110101000010010101010011110001010101001000111101110110000011110110011110011111011100110100111101110101010001110101010100110111010001010001011101010110100101110101001011010001010000101111101000000101010001111110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000100000000;
neuron_parameter[17] <= 368'b10010000000000000110111000010111101010010101011010101010010101110010100000101011100011001010101110000110101011111010010010101001101000011010100010100101011011010010100111010101101100010101000110101000010100011010101010101000101010101010101111111111100100000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000100010000;
neuron_parameter[18] <= 368'b00101010101011001110101110101011001111010100001000110101010100110001000010000010101000001010101110100010001010110011101101001011100110110100011001010010010001101101101100000011010100010100001010000101010110100110100111011010001010101010100000000010111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000100100000;
neuron_parameter[19] <= 368'b00010010101111010111011010101011100000000010101110000100110110111000010010010110100001100000001010100110000101110001001010110111100100101011001110010000101100101010010110010010001010100100001010101010010010111010101000101011101010101010100110100000110101010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000100110000;
neuron_parameter[20] <= 368'b00101010101011001010101010101000101010110101001000101001010100110000101100001111100010001010101010000010100010101001001011000011100100100101001010010101010100101000010100010010110100111001001010101001010000010010101001101000001010101010110000001100111101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000101000000;
neuron_parameter[21] <= 368'b01111010101000010010101010101000011011001010101111100100001010110110000000101011111100110010101110101001101010101010101010001010000110100010111100001001001010101010100100100011001010010010111010101000001010110010110000101000101000010010100010000011011100110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000101010000;
neuron_parameter[22] <= 368'b11001010101011010110110110101010100101011010111001010100100011000101011011010111010101100101010001010110100101100101011010110111010101001011011010101000100100101000101101010111101000110001010100101101010101010011010101010001011011010100000000010111110011010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000101100000;
neuron_parameter[23] <= 368'b10001010101010010010010000010010001011010100010110100100101101010011010010100101101101001010110010010010101010000000101101001010101011110010001010100100101011101010000100001111101001010110001010101011010001101010101011010011101010101010101100100010111011110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000101110000;
neuron_parameter[24] <= 368'b11101010101011110110101010000011000001011010001100001010100110100000100010101010101010001010101110101000001010101011010101011010100101011100001010110000110010101000001010001100110100101000101110001010100010101000101010101001001000101010101001111100100011000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001000110000000;
neuron_parameter[25] <= 368'b10001010101010001010100010101001001010101010101110101100100010101010100101010011101010000101001110101000000000111010101010010011101010101000101011000001000000101101010100101011110100101010101101001010101010111000101010101001001010101010010011101010100000110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000110010000;
neuron_parameter[26] <= 368'b01101010101000000110101010101011001011110010101100001011001010100010100000101011100100000000101011010001010100100000001101010010010100100101011111001001110101101001100101010110100110110100001010001010101011011001101010001101010101101001011000101100011001100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000110100000;
neuron_parameter[27] <= 368'b01110100000101001010110000000100101010101011011000101010010010100010101101001011101010010010101110000001000010100010110010101000101011001010110010101001111001010010110110110101101100011001010110101000100101010010101010101011011010101010111000111110011101000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000110110000;
neuron_parameter[28] <= 368'b10101010101011111110100000101010100101010010101000100110001010100001011000011011100100100000101110111010010010111011001001000011110100000101011001010010010101101001101011010010011101011101111011111100011010100110101001101001101010101010111000010110100101100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000111000000;
neuron_parameter[29] <= 368'b11100001010111110001000001010011100000101101011100001000100100111100000010011011100000111101001110100101010100100011000101000111100010010010101110100001101000101010100110101011101001010111001010100101010010100010101010101011101010101010111000000000100111110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001000111010000;
neuron_parameter[30] <= 368'b10000010101010000010101010101010100010100101001110101000001000100010100000001111101010001100111010100100110010111011011001000011101101100110101010111110011010101010110110101010001000001010101010111000001010111011011110101001001010100010011100001100101010110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001000111100000;
neuron_parameter[31] <= 368'b00101010101000010010101110101011111100010010001110010101101011100101010001101011110100100110101100101010011010111010100100001001001110010000111011101001101011101010100100011111001000001001011110110010010100111011000101001011101000110010100010011011111000110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001000111110000;
neuron_parameter[32] <= 368'b10101010101001010110101010100010100010110101011010001011010101111110100100010101010010010100010101101101011010100110100101101010001000000110101110100001001010101000000100101011001000010010011010100001101010101010000000101011111010001010010100010011101000110000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001001000000000;
neuron_parameter[33] <= 368'b11001010101010100110001101010110101101110010010010110101011010001001001100101100100000111010110010000001101011000011100100101010101011011100101010100101000000101010010110010111101000011001011010101011110100100010110101010011001011010110111101000110111110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001000010000;
neuron_parameter[34] <= 368'b11001010101011010100101010101001101100101010101010110010101010110011100101100000101101010110101110010101000110110001010000011001110101010101011110101100000001111010101000010010101010101001001111001010010110110100001000101001111010111010111111101100111100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001000100000;
neuron_parameter[35] <= 368'b00001010101010110000111110101110110001110110111101110100010010101101010011100011110101001011101010010110100010101010101001001110101010110101101011101001011000100110110100100110110011011001001001001001110110100100100100101000001011101010110110011100110111010000000000000000000000000011111111110000000011111111110000000110000000000000000000000000000000000001001000110000;
neuron_parameter[36] <= 368'b00101010101000011110101010101010101010101010101010111101010010110011000101010011110101010101001011000000100000101000100000000011100010010010001110001000101010111010101010101011101010101010101111000101010101011001010101010111010101010101011000101110011111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001001000000;
neuron_parameter[37] <= 368'b11110100010100001011110101001010001010100000101011101000011010100010100000101010101010010010101010001000100100111000100010001000101010101010100100101000101010010010110101010101001010010101000010101010010101011011101010101011001010101010101110000100111001000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001001010000;
neuron_parameter[38] <= 368'b10001010101011011010101010101011101010110111101000100010110110110010001010011010100110001101001111100010110100111011100100101010110101010010101001000011011010101000001001101011011001100110101011101001001010110010100110101010101010101010100111011000100111100000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001001001100000;
neuron_parameter[39] <= 368'b01010110010010111101010001011010110101101001011101010000101101110001010010101011101010101001001110101000110101110011010101010110101100010101011110001001000001101010100010100011101001011010001010100101101010000010101010101011001010101010101010111100100110110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001001110000;
neuron_parameter[40] <= 368'b10101010101011001010101010101010101010000100101110101000010010100010100010001010101000101000101000100110110010111011001010001010101100101000101100110010110010101011011000001011101001000110101010101001001010011011010000101011101010101010110010101000111100000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001010000000;
neuron_parameter[41] <= 368'b11011010101000100010101010101001011010100110001100101010000010101100001001001011111100100110101110111010011110101000101110111001100110111010111110101001101011101010110110101110101000111010111110110010101010001001010110101010101000011010101011001000000011100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001010010000;
neuron_parameter[42] <= 368'b01001010101011111010111010100000010101001001011101010010111001001101001001001010010110110101101101011011010100101100101100010110010110101011101111010100101101101001010010010111101101001001010110110010010100111010101001010001001010010100001011001111100010110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001010100000;
neuron_parameter[43] <= 368'b01001010101011101110000101011001001010100100010110110000010101011011011010010111101000001011010010010011001011001010000100101010101010010010101010001001001011001000110100101111100101011011010010010100101010101010101010001101101010010110111111111000111100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001010110000;
neuron_parameter[44] <= 368'b00101010101011101100101010101011111010110100101010001010010010100010101100101010101100110000001110111011011010101001101110011011100110011101101010111110111010101001111001101011110100100110101110011010011011100101001010101000101010101010110010110000101110000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001001011000000;
neuron_parameter[45] <= 368'b11101010101010001001010111001100000101000101101000011000010100110010000010100110101100101010111110111010101010110010001001001011101010100101111011101010010101100100101011001010110101010100101101010000111010101110111011101001001000101010101110001100101100010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001011010000;
neuron_parameter[46] <= 368'b00101010101010110010101010101010001001001010101000110101010010100010101101001011110001010101001011010001010100111100100010000010110010010000101010001001001010101010101000101010001010101010101111101010100101100001010101010111010101010101010000100100001100000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001011100000;
neuron_parameter[47] <= 368'b10011101000101011011100111101100001010011010011000101001101010101010100110101010101000011010101010110100101100111001001010001101100100001000010010100000010000010011000101010000100110101001000110101010101100010010101010101001011010101010111100010000111000110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001011110000;
neuron_parameter[48] <= 368'b01001010101010101010101110011001100111000001101100010010010000100000101001001011100010110100101110001001010110110100100101101010101110010101001101010001010011101001010010101010010101001010101110101100011100101000000101111010101010101010100000111111101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001100000000;
neuron_parameter[49] <= 368'b01000110101010100011000010101011100010101010101010001010000010111010000101110011101000010101011110100101010101110001010101000010100101010100011010010101000010101001101010101011100010100110101010101011010010100010101100101010011010101010000110111011111010100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001100010000;
neuron_parameter[50] <= 368'b00001010101011100010101010101010001010100011101100101010101100110010101001011010101010001011111000110100111110111011011011011010101101100111101000111110011010101011110000101011001100001010101110101001101010100010011110101000001010100010101001100010101111110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001001100100000;
neuron_parameter[51] <= 368'b10101010100111101110101010101000111011100100101110101010000010100101011001001010110100100010101010111010101010111000101110101000100110111010111010001001101010101010100110000010001010001010101010101101101010110010110010101000001000010010111000100100100100110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001100110000;
neuron_parameter[52] <= 368'b10001010101010011010101010101011001110101010101011110010101011001010101010100100010000001011010101010101000101111101010101010110010000100100101010110010101010101001001010101010111100001010101110100100001010001011000101001000011010001100101111011111101100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001101000000;
neuron_parameter[53] <= 368'b01101010101011011010101001010111001010000101010000101000000101010010010010100100101001001010100010101000001010010010101001001011101010000010111010110100101001001010010010000101001000000000101100100100010110111010101011000111001010101010111111110100010111010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001001101010000;
neuron_parameter[54] <= 368'b01101010101011001100101010000000000100010100101000010000111010101010100010101000101010001010101110000001010110100001100101000110111111001101001010101000110010001010100000100001110100101000011010010000100101110100101010101010001010101010100101010010110001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001101100000;
neuron_parameter[55] <= 368'b00101010101010000001100011001100101010001101011000110000010100111001001011010010100100101001011110000010100101101001000001010111110110100101011011011010010010100101001000101010110101100000001000010101100010111001010110101011001111101010111001110011100010100000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001001101110000;
neuron_parameter[56] <= 368'b10001010101001010010101010101011101010101010101000100100001010110100001001000010110000111101101111000110000000101001000110000011100100001101101010010000110110111010101001101011101010100100101010101001001010010010100101100111010011010101001011011100010000100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001001110000000;
neuron_parameter[57] <= 368'b10110000001101101010010110100101001010001010101010111010010101100010101001011011100111010110111110010100100101101101011010110100100101001011010010101001100101010011010110010101101011000101010110101011110110011010101010101000001010101010100011001101101111110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001110010000;
neuron_parameter[58] <= 368'b00001010101011000110100001101011001010010100011100001010100100111001101011010011100010101101101110001010010000111110100100101011110100000000101101000110010110101001001000011110010000111111011110010000011011101001011000101010101011101010101000111010100111000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001001110100000;
neuron_parameter[59] <= 368'b11000111110110100011010010110111100100001010101000111010101011100110100010101011101010001001101010101000010011101010010000010110101101000101011110110100110101101010110011001011101001001110101010100010011010110010101010101000101010101010100111111110111010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001110110000;
neuron_parameter[60] <= 368'b01001010101010011110101010101001001000010001101010101000000100101000101001010111100100101011011000010010101101111000101010110110110110101000001010001010111010101001001000100111100111000000001010000010010010011000001000101010111010101010101100001100101011110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001111000000;
neuron_parameter[61] <= 368'b01111010101111101110101010100001001000001011001101100100100101101000010110011011101000011000101110101010101010101010101110101011101010101011011010101010100111101010011001001011101100100100111000010010010010101001101100011010001000010010110001000000111111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001001111010000;
neuron_parameter[62] <= 368'b10001010101001010110101010101000001010101010100111001010101011101101000011101100010101011001010001010001000001011101100101000011010011010010101010101001100000101010101100000011011010101010100010101010101000110110101011010000101010010100011001110001101011100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001001111100000;
neuron_parameter[63] <= 368'b00001010101011010110101101010010101000000100010100100001010011000001000101000010100010000110110110000001001011010000100100101111001010010010101110101011001000101001010100100001100101010011000010100001110101110010111000010011101010010010100011000000101100100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001001111110000;
neuron_parameter[64] <= 368'b11101010101010010000110010101010101101011010101110110100101010111011010000101001100101100110101011010101001110111111010101001011101011000101011110101000010100101010101001010011100010100101001110001000000100010101101100001000101010101010111100100000100100010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010000000000;
neuron_parameter[65] <= 368'b01101010101000001101011001011010110010101101011100000010010101110010000011010101101001010111011110000000001101110001010011010011110100101101011011010010100100100101001011010011010101100100101000010100100010101001010010111010001111101010100010010100100001000000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001010000010000;
neuron_parameter[66] <= 368'b11100010100111010110101010101001101010000000100010101000110010100010100000001010101011001100101010101010010010100010101001001010101010100110101110101011001010101010100010101010100100001011101011000110101010111001011010101001100101110101001011000000001100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010000100000;
neuron_parameter[67] <= 368'b11010001010100100111010101000001001000010010101100111010101010110010101010101010101010000110101010111001010111100001100010010100100001001001010010010100100100010001001111001101001101110100010100101010110101011010101010101010001010101010110111101101100001010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010000110000;
neuron_parameter[68] <= 368'b11001010101010011010101010101001001001010100101110010101010100100001010001010011100000100101001010101010001010111011101110101011100100001010011101100000100000101000000001010011000101010101101010110101010000101110010100011001001011101010101101001101100001000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010001000000;
neuron_parameter[69] <= 368'b01000100101110101101011110010001000101100110111110001000101011110100001010101110110000101010101010110010101011101011001010100111100100010111011010010101001101101010110011010010101010110100101000101001010010100010101000101010011010101010111101010000110110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010001010000;
neuron_parameter[70] <= 368'b11001010101010011010101010101010001110110010001000101000110100110000000101010110100001000101011110000010100101111101001010101011110000100010001010000101001010101000000100101011101011011100001110000101010000010000100101001011101010101010110110000001110000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010001100000;
neuron_parameter[71] <= 368'b10001010101101111110101000101000101111011010101101110000001010100001010100101011101100010010101110101010101010101010101010001011001100100001101110011010011110101010101101100011101010110010101100101001011010110010101101001010101010010010110001001111001101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010001110000;
neuron_parameter[72] <= 368'b10101010101001011010101010101001101010101010101101001010101100101001100010110010010101001001011001010101010101111100000001000110010000100000101110100010101010101010001010101010111000100010100010101100001011010110100001010010111010001100111010100001111100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010010000000;
neuron_parameter[73] <= 368'b01001010101010101011010101000110101101010110000110111100011010000000100100111010101011001010111110010100101001000001010010010111101101100101001100110100100101011011010010010111001001001101010010101010010101011010010101010100101010001110110000000100101101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010010010000;
neuron_parameter[74] <= 368'b10001010101011010110001010100000100101100001101000001110001010101010101000101010101010100010101110101001010100100001010100010010101001111101011110101110110101111010001010000000100010101000001110000010111001111101001010011010101010101010110111100100101100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010010100000;
neuron_parameter[75] <= 368'b00001010101011101100011101101001110011010000101110010011001000111000001100101011100010110010001110001001001010111010101101000010101010010100011011101011010100100101101001010010110100110100101001010011111110101011101010101000001011101010111111101101110101010000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001010010110000;
neuron_parameter[76] <= 368'b10101010101000111010101010101001101011111010101010111001001010110000100110101011101010010100101111010001010110100101001101011010010100110001101111111010010110101010101101001011100110100010101011000010101010011101001010100001010101100001001111010010000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010011000000;
neuron_parameter[77] <= 368'b11110010000100011011000001011101001010000011011111100100000000101010000000101010101000001010111000110010101101111110001010000000101001101101000110010110010001010001010000100001000010101010110110001010101010010010101010101000111010101010000001110100111111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010011010000;
neuron_parameter[78] <= 368'b01000010101011110110100001001000001010100100101000111010000110100011100110011010101010111100101110101010011000101000000000101011100100101000001001011110110110101100101000101010010100011010101011000100101010000110111010101001101011101010011010000100000011000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001010011100000;
neuron_parameter[79] <= 368'b00101101010110111111010101010110100100000101001110110000011010100010000001100011101000000110101010101010001010111010100010101110101000001000011110100100100100101010010101010010101101010100101110110110111010100010101010101001001010101010101110110010101111100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010011110000;
neuron_parameter[80] <= 368'b01001010101010011110101010101010101010110100101100101000010010101010001011001010101100001001101100100110100010101011001010001110101001101000101110110110100010101010010010001011001001001110101110101101011010110011110100101000001010101010010111101110100011110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010100000000;
neuron_parameter[81] <= 368'b10111010101010011010101010101000011000001010001011110100110101110101000001010010100000110000101010101011101010110000100110101000101010010111011110011001001011101010100100111110100100111011011110000010101110101001001001001010101000000010110110010010101100010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010100010000;
neuron_parameter[82] <= 368'b01101010101011110110111010100010011100101101011111001010010100101001101101010011010010010100010101101011011001101010000100101011011100111010101011110100101000101011010110101010101100111110000110111000000010100010101000000001001010011010110101110011111001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010100100000;
neuron_parameter[83] <= 368'b01001010101010101010101010010101101000001100000110101010010001011000100101010101001001001011010010110010101001010001001010000011101010000100001000101101001010101010010010101100101001001010111010100100000100101010000101010100101010000010100001011110000111000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001010100110000;
neuron_parameter[84] <= 368'b01001010101011111100101010000001100011010000101010001010000010100010100010101010101010100010101010101001001010100010010101001111100001010101101110110100000010101000101000111000100000101010101110011010101111100000101010101001101000101010111001100110101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010101000000;
neuron_parameter[85] <= 368'b00101010101001011101010101111001010101010010101101000001011000101000000101101000111010110110101110000001001010100000110100101011101001010110011001001001010100100110101101000011110010010010011000001010000100001100101010100000001010001010110001101100111000110000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001010101010000;
neuron_parameter[86] <= 368'b00001010101011000010101010101011101010101010101110110001010110110001110101001010110100000000001010000010000000101001000101000011100100000101011110010010110001111011001010100011101100101010101011010100101001011001010100000010100101010101001000111010000001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010101100000;
neuron_parameter[87] <= 368'b01010101010100100011010110011111101010011010001011101001101010101010100110101011101000001010111000000000101010111001001010000001101000101000000000000000010000010001100101010101000010000001000110111010101011011010101010101001001010101010100000010010011101110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010101110000;
neuron_parameter[88] <= 368'b00001010101011100110000100101011001010010110101011101110100010100010110011001010101010010110101010101001001010110000101100101011101001100101101000110110110010101110000011001010001000100010001111100100101010110110000010101000101011101010110110011110100110000000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001010110000000;
neuron_parameter[89] <= 368'b10000011110110000001111101001010000110100110101100111010001010110101100100101011111010001000101100101000010001101010010100101100101101101000111110110010110010101010000000101010101001011010101100100000101010011010101010101000001010101010111110111100111101100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001010110010000;
neuron_parameter[90] <= 368'b11101010101010100010101010101011001010010100101110101001010100100001001001000011100100101000001111000010100000101001001011000010100100100101001110100101010010101010000110110010101010101000001110110101010000100000110110101000001010101010111101011110101000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010110100000;
neuron_parameter[91] <= 368'b11101010101101100010101000101001111011001001000100101000101000101100101011010010111010100000101010101011000010100010101100101011000110110010111110101101101011111011100010101111101001101010111010011010101010111011011110001001011010011010100010100000000000000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010110110000;
neuron_parameter[92] <= 368'b10101010101010001010010110101000110000000000001111010010010000100101100001001011010000000100101101011010001010110010100010101011110011001010101011101000100001101010100101010011101010100101010000101010010000100110101011010001010010101000101100111011110111000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010111000000;
neuron_parameter[93] <= 368'b10101010101010001110101000110010101101001101010010010101100101000000010010010101100100001011011010000010111011001010101100100110101010010010101110100001011011101001000101101111101100100110001010110001010011100010110100100000001010001010100001101010111110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010111010000;
neuron_parameter[94] <= 368'b10101010101011001010101010101011111000111100101010010010001010100011001010101010101000000010101010100011111000111010011000000110100001101110101110100110011010101011011001101011110100100110111111010010011111110101001011101000001010101010110011110010100101010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001010111100000;
neuron_parameter[95] <= 368'b11001010101011111001110101011110110101010000011101010101010110110001000100100010100101001010011010000010101010100100001010010111101010101001011011101010010100100101101101001011110100110010101101010001010100100101001001100001101001001010101110000000100001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010111110000;
neuron_parameter[96] <= 368'b00101010101010101110101010101011101000101010101010110001000110101011000101000010110000100100101110000101010110110001000100010011110110011101101010100010100011101010101010001010101110101010111011010000101001101001010010000110100101010101011101110100000111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011000000000;
neuron_parameter[97] <= 368'b01110000000100010111000001011111101000000010101111100000001010110010100000101011101000001010111100010000101011110100001010000001101000001001010100110110010001010000010001010101000010101011000110000010101011011010101010101000001010101010100110110110110101100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011000010000;
neuron_parameter[98] <= 368'b01101010101000110110010110011010101110001000101100111010101010110000000001000110100000010101001111010001010100100110010101010011110101010101101101010101010100111101010001000110000000101010111110101010101010111010000000101000101010101010110001010100111001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011000100000;
neuron_parameter[99] <= 368'b01000101010110111001010101001011001010101000101000001010101010100000101000101011101010001010101000101000010010110010100101001011101011010001101110100010110110101010001101101010101000010010101100100000101010000010101010101010001010101010010110010000110000000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011000110000;
neuron_parameter[100] <= 368'b01001010101011101110101010101010001010101101101110101010100100101010101001001111101011001101101110110110110110111101011001011010110100100101101110000110011010101010000100101010000000000010101110101000101010011010000010101000001010101010110101001010101001100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011001000000;
neuron_parameter[101] <= 368'b00101010101001111110101010111001001101101001001001000100010100101001100101010010101000011000101010101000101010101010100000001010101010010010011110011011001010101010100100101011000101001010011110010000101000110001010100111001101000000010100000111110100100110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011001010000;
neuron_parameter[102] <= 368'b00001010101011100010000100101001010101010100001111010100001101011101010001000110011010000000111100101010000010111010101010101010101000101010101110010010101000101001011000001111100101000011111010110100000110100111010001001000110011010101000101101101110001100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011001100000;
neuron_parameter[103] <= 368'b10001010101010011010011101010110101011011001010110101010101101000010110100000101001101011010010110100010101011011010011100101011101011111010101100100101101011101011010110010100101000110101011010101111000101110010010101110111001010001010100111010010111000110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011001110000;
neuron_parameter[104] <= 368'b11001010101010011100101010100011101010101010101000101010101010100010100000001010100001010101001111000001100100110001010001010110110100000101011010010001010101101000000010000011100000101010101110101010101000101100000000000000101010101010110111101110101110100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011010000000;
neuron_parameter[105] <= 368'b11001010101010110100000100011101110010000101101001010100101000100101010010101011100110101010101110001010010010110000101001010011111010100101011111101010110100100101001011000011110101001101001100000000110010101101100001100010001000101010101111011000111111110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011010010000;
neuron_parameter[106] <= 368'b00101010101011011110101010101010101010101010101010101010001010110010100001101011101001000110101010110000110010101011010011001011101101000110101010100010011010111010101000101010101010110010101010101000001000000010010000101010010101010111010100101110001100000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011010100000;
neuron_parameter[107] <= 368'b11010101011101000110000101010101101010000101011110101000101010100010100010101010101000101010111110110101101000111000000111101101100111011110110110110101010010010011000101000000001011010000100110101001100000011010101010101001101010101010100100111000100110100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011010110000;
neuron_parameter[108] <= 368'b00001010101010010110101010101010101101010100101000110101010101101001010010010111101001001001001110100010101000110010101000100011100100101001011000010010010100111101001001000010010101010100101010000101010110110110010111001001001010101010100001001000100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011000000;
neuron_parameter[109] <= 368'b11100101001011011110110111011000011011001000101110001010001010110000101000101011111010001010101010101000111010100010100101001011101011010101101111101101100110101010111011001011101010010010101000101000101010101010101010101000001010101010010111001100110111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011011010000;
neuron_parameter[110] <= 368'b10101010101011101010101010101010101011010001011000101001010101101000001101010111100000000000001011000010100000111010001010101010100000101010001010100101010010101010010100100011100001010000001110010101010100100000110100001010101010101010100110111100100110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011011100000;
neuron_parameter[111] <= 368'b01101010100001011010101000101010111010001100000100101010101000101100101011010011111000100100101110101010010010101000101100101000100110111010111010100101101011101010100010101110101001101010111010010010101010011010011110101001001010011010101100111010000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011110000;
neuron_parameter[112] <= 368'b00001010101000011010100010101000101100000010101001010100010101100101010101010111010100011001011000101010101001100010001010101110101000001010101110100010101011101000000010100010100100010000001010100101010101100010010101010001111010010000101111101111110000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011100000000;
neuron_parameter[113] <= 368'b01001010101010111010000101010100001001000001100010110110101101000001011010000111100100101010110010010010000010000011000000001011001010000010101010100010001000101010100000000111101010110110001010101010100101101010101010111101001010101110111010011111111110110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011100010000;
neuron_parameter[114] <= 368'b10101010101010100000100000101010000010001011101111000010100010110010101010101010101010101010101010101010001010110010010101001110100101010111101110100110110010101010011011001101110101101100101010010010110111111000101010100001101000101010100111110110111001010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011100100000;
neuron_parameter[115] <= 368'b11001010101010001101000000011001010101000000011001010000010101100111000000001111100100001010011110100000101010100010000100101110101010010000111010101010101110100010101000101011110101010110101001010100011010001101011010101010001001001010010011110100101100000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011100110000;
neuron_parameter[116] <= 368'b11001010101011110110101010101011001011111010100110011000101010110001100000001010100101010101001010010100010100111000001001010010100100110100011010010011010101101001100101100010100110111010101011001010101011100000001010001111010101010001110111110110001010100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011101000000;
neuron_parameter[117] <= 368'b10011000000100110010010000011101001000001010011111100000101000111110100010101011101000001010101010001000101000111001001010000001100001001101000010010100010001010001000001000100000110000010010110111010101011000010101010101001110010101010101000110001101010010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011101010000;
neuron_parameter[118] <= 368'b10101010101011000010101000111011001010100101101001110010011100110001101010110011100010101001001101001010010100111100100001101001100101000000101001011010101010101001101100101011010000011010101111111100011010000010100000101001001010101010001001111100100110000000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001011101100000;
neuron_parameter[119] <= 368'b11000001001110110100110101101000011010001010101101101000101010101000100010101011111010001100101100101000110010111010100010101011101011010001101110100100110010101010110011001010101010010110101100101001001010111010101010101000001010101010110010101110100111010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011101110000;
neuron_parameter[120] <= 368'b10101010101011110010101010101011101001001010101000010100101000101010010010000011100101001101011010000100110101101000011001010011100011101000001010000010101001101001010001011011100101010110101010010100001010101011101001001010101010101010101001101101101100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011110000000;
neuron_parameter[121] <= 368'b01101010101010111110101010011010001000100101001101000011000101110000000110010011111010001010101110101001001010110010100100101010000010010010111010011100011010101011101000101011001101010010101010010101001000001010010010101001001000000010110010100100111111000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011110010000;
neuron_parameter[122] <= 368'b01101010101010011010010110101000010101000001001011010101010101000101000101100010010010100100101100101010001010111010101010101010101010101010101110001000100001101001000100000110100100010111110010110000010001100110101000000000010010101001000101111101110000010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011110100000;
neuron_parameter[123] <= 368'b01001010101011011110001011010000001010100100000010100011000011000001010000010010100100001010100110010110101010001001000010011010101010110100001000101001001011101010110110101101101010001001010110101001010001111010101101000101101010101110100110111111101111110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001011110110000;
neuron_parameter[124] <= 368'b10101010101000101010101010101011000001101010101001100100101010101010000010101000101010011000101010100000000110111011000011000111101010001101001010101000000010001010110010000000001001001000011100100100100001111011010010101000101010101010100010011010101100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011111000000;
neuron_parameter[125] <= 368'b11101010101010001011100000101001001000001001011100010111100101111001000010010000100101001001011110000110111101110011101001010111111110100100011111011011001000101101011010010011110101100000101001010101101010100101010010101011001011101010111000000001110011000000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001011111010000;
neuron_parameter[126] <= 368'b10001010101010101110101010101001001010001010101110100101010110100011010101010010111001010000101110000000100000111100100001100011100001000000001110100110001010111010001010100110101101111000001011010101010101110001010101010100010101010101011000010010000100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011111100000;
neuron_parameter[127] <= 368'b10110010001001111111000111111100001010011000001001100011001010111010101000101010101000111010101010101010101011100001001010000100100010101001010110000111010000010001010100000000001000101001010110111010101011011010101010101000011010101010101001110100000100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011111110000;
neuron_parameter[128] <= 368'b01101010101011111010110010101011100101000000001110110000100000110000001011010011101010100101001110101010010010101010100100101010110001010010001101000100000100101001011010000011001101100000101010110001010010110101001000101000101010101010101111011010111000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100000000000;
neuron_parameter[129] <= 368'b10100111111110001001011110010100100100101001101000001010001010111000000000101011101000100100101110100010000100110010011101010110101101101011011110110110101100101010011100100110101001001000001010100100100010100010101010101001001010101010101011111010110011010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001100000010000;
neuron_parameter[130] <= 368'b00101010101000000010101010101010101011010101101110011011010010110010101001001010100010100100101010001010110010101001001011010010100100101101011110010010000101111000010101010011100101010010101010100110101010101000100011101001001010101010111101110110110000110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100000100000;
neuron_parameter[131] <= 368'b11011010101001010100101000101001001001011010100011100000001010100000010100111010101110011010101010101001101010110010101010001011101110100100111110111010011111101010101101101111001010110010111010101011011010110010101100001011001010010010111111010101101110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100000110000;
neuron_parameter[132] <= 368'b00001010101011100110101010100011001110101101001010001010010100001100101101000000010010010101010101000101001001111110101100101010011010010010101010100001101000101000010110101110100111011010110010001100100011111010001000000001101010111010000110011001101100100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100001000000;
neuron_parameter[133] <= 368'b11101010101011010110001100011001001000010100010100000000110101101000000011010110100000101101001010001010011111000010100100101111101000010110101100100101011011101010100101101010000001010010101010010100001011101011001000100011011010001010111010010010101100110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100001010000;
neuron_parameter[134] <= 368'b11101010101011011010001010101001000000001010101011010000101010101000000010101010001010001010101010101000001000110011010100100110101100000001001010101100100110001010010010010011001001101001011010110110100101111001011010001001101000101010110100100100100000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100001100000;
neuron_parameter[135] <= 368'b11101010101001111000100101001111000010000101011100010011010101101001001011010100100010001001011010101000000101110000010011010111111101101101011011010110100100110101011011001010110101100000101101010101000010100101010110101011001101001010101100010011110100100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100001110000;
neuron_parameter[136] <= 368'b00001010101010110110101010101010001010101010101000101010100110111010000100011011111011010111101111111111011100110001000001100011110100010001001110000000001010101010001010100010101010101001001111101010100101111100011000010110010101011101000110110100000011100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100010000000;
neuron_parameter[137] <= 368'b00010101010101001110010101010111101011010101001000101001001010111010100010101011101010100010101110101001011010111011001111111001101100001101110010110100100110010001010011010100001100111101000110101010010101010010101010101000101010101010111111011001111001000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100010010000;
neuron_parameter[138] <= 368'b10101010101011101010101111101011001101010100101000110101001000111011000010111010100010000101101010001001010110100100101101101010110010100010111101011011010101101100001101010111010010010001011010010101001010101001100001101010001010101010110010110111100100000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100010100000;
neuron_parameter[139] <= 368'b00100101011110100001110101010101011010101001101110101010001011101000101000101011111010110110101100101111000111100010110110111011101101001101101010100110010010101010001101101010100110010010101110101000101010010010101010101011101010101010100101111110110000110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100010110000;
neuron_parameter[140] <= 368'b10101010101010000110101010111001001010000010101010000001001010110011000101101010100010001100101101000000110011110110111011101110100001101010011010101110011000101010110001001010101010010001001010101010000010100010101110001011111010101010100101110110010110100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001100011000000;
neuron_parameter[141] <= 368'b10011010101001000010101010101001101100101000001111000110010100110101100100010010101010011010101110101001001010110000100100001001101010010010011010011001001010101010100100111111100100101000111010010000101000100001010110101001101000000010101000111100011001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100011010000;
neuron_parameter[142] <= 368'b11001010101011001010101010101011101010101010101111010010000001111101010011000111010100000101011001010000010101011100100101000110011010000010101010101000101010101010100010001010101010001010100100101000010001011010100101000011011010111100011011010011110001010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100011100000;
neuron_parameter[143] <= 368'b00111010101011010010101010101001101010101010110010101000010110111010100101010100001011000011010010100110101011000011110010101010101010000000001100100101000010101001000010101011001101101010101110110000101010100010110101011100101010110010110010101101100010000000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001100011110000;
neuron_parameter[144] <= 368'b00001010101010101000101011000011001010100100101110000000010100110010000010010110101000011001011010101000110101111010000001010111101100000100001010110000110010101001000000101011010101001010001001010100100010111101000101101011101110101010100000111110100100100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100100000000;
neuron_parameter[145] <= 368'b00001010101011110100110100101010100000000000101000010010101010101001101000011010100010010100001010101010001000100010101010010011101010100101001111010001010100101101010110111010110100101011001100101010101100100010101010101011001010101010110010100010101101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100100010000;
neuron_parameter[146] <= 368'b11101010101011111010101010101000101010101010100110101001001010101000110101101011101011010110101110000000011000100001000100100011110100011000001110010000101000101000001010010010101010101101101010101010000001111010100100010110000111010101001100110000001110110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100100100000;
neuron_parameter[147] <= 368'b01110001010000000010001001010110001010101001011100100000110000101010101000101011101000100010101000100010101010100000000010100001101101001001010110010100000101010011011000010001100001001010100100101010010011000010101010101001101010101010000001001110101001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100100110000;
neuron_parameter[148] <= 368'b11001010101010000010101010011010000010000011101000110010011100100001001010110010100110101001001011000010110100110101000011001011100000010010101100011001011000101001000001011011010001001000101011111000011010100110100000101010001010101010111100010010111100100000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001100101000000;
neuron_parameter[149] <= 368'b11010110001111111001000001011010010010001011101000000000111010100010001011101011100001001100001010100000110001100001000001010010100101010101001110010111010010101001001001101011110110110100101010101011010010101010101100101001111010101010100110000010100101110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100101010000;
neuron_parameter[150] <= 368'b00001010101011001110101000101010001001010101011100110110010000111000100101101010101010010100101110100000110100110000001010010110100100101000011000000010100101101001010101011010100101010100101010000000101010001010101011001010001010101010101110110010111011010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100101100000;
neuron_parameter[151] <= 368'b00111010100100100110101010101011011010100001100001110010010011111101011001001011110000100010101110101010101110101000100010111011000110011011011010001001100111101010110110000111001001011010111100100001101010000011010110101000101000010010110110011001000000100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100101110000;
neuron_parameter[152] <= 368'b00101010101010110010110010101010011101101010101101010010111000100101010001001011010110000101101101011010010110001101101000101010010111001010101011101110101100101010110000010111001010000001111010101000010100100010110001010011011010100100110010101101101111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100110000000;
neuron_parameter[153] <= 368'b00101010101011110110101001010101001010101101010000100100110101001010010011000110100000001100100010001010011001000010000100101011101000010010001100100101001011101011010110100111101001001110010010101000110011111010111101000110001010010010100011110001111111110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100110010000;
neuron_parameter[154] <= 368'b01101010101011001010101010101010101010111100101100100000101010111010101100100101101101010010001010010101110110111110100010011010101010000111101010101110011010101010001001101010100000100110101011011010001111101100101100101001101010101010111010100100111000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100110100000;
neuron_parameter[155] <= 368'b00101010101010011010101010101011111000101010101011000000010010101101101101010011100010010000011010010010101001101000001010101011101101010110001011010001001010101100101010111010101010101111001000000101000100100001010100111011101000001010111010000100100011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100110110000;
neuron_parameter[156] <= 368'b11101010101011001110101010101000101011001010100000000010001010101000010001001011100000010101001110000100010100100000001001010011100100101001011010010010010001101001101010001010000100101010101111010010101010110011000010001101000101010101010001001000001010000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100111000000;
neuron_parameter[157] <= 368'b01110101000001011010100101010101001010100001011101101010010011110010101010101011101010100010111100111110101001111101011010000100101101001010010110100101110011010001010000000100001001010100110110101010101010001011101010101001011010101010010101001100110010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001100111010000;
neuron_parameter[158] <= 368'b01101010101010111010101010101001101110000001011000110000110000100001001011001011101010100100001010101010010010100100000001001010110100010010101001010101000011101001010010001111000101101010101110010110000010101010000100101001001011101010110000011011101010110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001100111100000;
neuron_parameter[159] <= 368'b10000110010111101111010000000011000100001010001110000000101010110000010010101010101001010010101010101001001001110010000100010110101101010001011110110001110101101001100010010111110011001010101110101101101010111010101010101001101010101010100010100110110011100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001100111110000;
neuron_parameter[160] <= 368'b00001010101010110110101011101000101010100000001110001011000000101001000001101011100010001000101010010100100100111000011011010110110100101101001010010010010110101001010101001010000010010010101010101010101000011010000001101010001010101010110100111110110100000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101000000000;
neuron_parameter[161] <= 368'b10011010101010101010101110101000111101001000101000010100100101110101001100111010110100110100101110101011001000111000100100101010001110010001011110101001001111101010110100110111100110001001011010001010010100101011000100001000001010100010111110011101110001110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001101000010000;
neuron_parameter[162] <= 368'b00001010101001110110101010101011001010101010101111011010100100111101010000110010010101010101001101000101010100100100000101000010011000100010101010100010101010101010001010001010101010010010100100101000100100111010100111010100001010110100101001111011111111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101000100000;
neuron_parameter[163] <= 368'b11101010101010001110010001010111001111000101010000111101100011011011100010110101100101001001010110010110000101000011011001110110101101100100011010110110100101001001101011000110001010100110010110000101010100101010010101110001101010001110100011010111111000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101000110000;
neuron_parameter[164] <= 368'b11101010101010010010100000101010000001100010101100010010001000101010010000100000101000011001011110010000101100100010000010010111101100001000001110101100110000101010011010001101101101101001011010010010110000101111010010101011001010101010110001010010111100010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001101001000000;
neuron_parameter[165] <= 368'b00001010101001011100000001011001010100010100001101010001010010110100100010100001110100001010001000010010101011110001001000101111101000101011001000101010110110100110101001000010110100010000101001010101001110101101010110011011101101001010101110011001101100010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101001010000;
neuron_parameter[166] <= 368'b10101010101011010010101010101011101010101010100010101001001010111000110001101011110000000111001110011010111000110001100011110001010110001011001110010010100100111000001010000110101010101000001010101000110101001010010001010100000011110101010001000010010010010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101001100000;
neuron_parameter[167] <= 368'b01010100000001101111000010011111001000001000011011100000100010111010100010001010101000001000101100110000101010100001000010000101101001001000010100010111010100010000010001010101100000101010010110101010101011001010101010101001010010101010100000110100001111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101001110000;
neuron_parameter[168] <= 368'b01101010101011001010101111001010100100010100011110101001010000100000101100101010100010000010101110100100101010110110010101001010100111010101011000001011010111101001100100101010010100010000001011000001011010110001100111001001001010101010101001111100111101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101010000000;
neuron_parameter[169] <= 368'b00100001010111001101011000010100000010101010101000011010001010110100101010101010111010000001101000101010010110111010001100010010101101001011011110111010010000101010001100101010101001011000101000100110101010011010101010101000101010101010010000100010100011100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001101010010000;
neuron_parameter[170] <= 368'b01101010101010101010101000101000101110010010101010000011001010100000000101001010101000000101011110100010100101110110001010010111110100101000001110010000001010101010000110100010100001010010001010110100100010010010001000001001001010101010111110111100101001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101010100000;
neuron_parameter[171] <= 368'b10101010101111100110101010001011011010001000000100101010101000110110101010101011111010101101101010101010010110110001100110101010000110111010111010100001101011101010010010101111101101101010111010010110101010111011001010101011001010101010000010001111110010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101010110000;
neuron_parameter[172] <= 368'b10101010101011000110000110101010010100000101101101010000010010001100000101011010010010100000101100101010100010100010101000001010101010101010101110101110101011101010010010100110101011011000011110101001010110001010100101010010011010100100001101011001111001100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001101011000000;
neuron_parameter[173] <= 368'b10001010101011000011010100010101001100100001010110000000100100011001000110110100100101011010010010010100101101001001011010010110101101101011011110110100101101001011010010110111101010010001011010101001010101101010010101010101101010101110100000000010111001100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001101011010000;
neuron_parameter[174] <= 368'b11101010101011000010100000001000111101010101101000110100101100101011010000100110101001000110011110101001011111111010110101010111101010001101001110100010100000101010101010001011101101010100001111010101001001101000000010101011001010101010100001110010111010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101011100000;
neuron_parameter[175] <= 368'b11001010101010011010100010101000011010101010101000101010010000110010101101010010101001001001011110100110101001100010000000100110101010010110101011010001011010101100001001101011110010101110101000100010101010110000011101101000001011101010001100011101111000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101011110000;
neuron_parameter[176] <= 368'b00101010100011000010101010101000001010001010100100000000011010111101001011001011100010101100101010110001110110101011001011001010101100001100101010101010010010111010101001101010101010000110101010100000001010110010010110101011010101010111000100110100011101010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001101100000000;
neuron_parameter[177] <= 368'b00110011000101010111010000010100001010101011001000101000101010111010101000001010101000010100001010100101000101110001011010110101101101001010010010110101001001010010110100000100101001011101100110100010100010010010101010101010101010101010101001111011100011000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001101100010000;
neuron_parameter[178] <= 368'b11101010101010000110110110101010101101001010101100110011101010100011001111101011101111011110101111100011111010101110101100101010100010111101001000100111110101111010011110110110001111111001101010100001100010100101011001101011101011101010111110010010100010100000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001101100100000;
neuron_parameter[179] <= 368'b01000101010110011101010101010000000100001101001000010000000110101100000010101011101000010010001110101000101010101010100010001111101001001001011010110110010101101001000101000010100100010100101010111001010010101010101010101011101010101010111011010000100100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101100110000;
neuron_parameter[180] <= 368'b01001010101011101010101010101011001011000010101010100100101000101010010000000110101001101100001000000010100100100001001010010110110100101001001100010010110100101001010001001010101110000100101010101011011000101010101001001010001010101010101010110100101000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101101000000;
neuron_parameter[181] <= 368'b10001010101110111010101010001010111010100100001100101010101000100110101000001010111010100100101010101010010110111000100110101010100110011010111010100101101011101010110010101110001101101010111110000000101010011000011010101001001010101010001101001000010010000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101101010000;
neuron_parameter[182] <= 368'b00101010101010100110010110101010110101011010111011010100100011110101010001010111010101101101010001010110110101011101110010010111010110001011001110101000110101101010101001010110101010010001011110100101010101110010010101010001111011010100000100011101100110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101101100000;
neuron_parameter[183] <= 368'b00101010101011100010010100100000001111011000110010101001001100111000100110110100100100011011010110000101100100001000010011001010101001010110101010010101001010011001010100100101101010110011011110100100100101101010101000010001001010101010101000100010111001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101101110000;
neuron_parameter[184] <= 368'b11101010101010001010101010101011010001001010101000100100101010111010000010100101101000011000001110100000110000110011000011011100101010001100001010101001001011001010100010101110101011001010011010101100101001100011110110101001101010101010110101110000110110000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101110000000;
neuron_parameter[185] <= 368'b10001010101011111010101011101000001010000100111000101000000101101010100000000010101011000001001010101100101000100010101000001011101010100110101011001000011010100101000101101011110100000010101101010010001010101100101010101001101001101010101000001010000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001101110010000;
neuron_parameter[186] <= 368'b11101010101000011110101010101000101010101010101000101000101010111000000100100010110110010010101011000011100000111001000110000011010101001000001010010100110110101010001011000011001010100100101010101010000000101010101101000100000011010101011111110100010001110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001101110100000;
neuron_parameter[187] <= 368'b11010101010101110110101101011000001010110101101011101011001010100010101100101010101010010010101110101000101010101101011010000000101010101010010010101000101011011010010100000101101101000100110110101100011010011011101010101001011010101010001100111001100110110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101110110000;
neuron_parameter[188] <= 368'b01101010101011010010101011011001101101010101101100110000010100100000001001000010101010100101001010101011001010110010101100101010110100010010011001010101101101101001010010010010011101000101101110000100010110100000111101011000001011101010100010000110100001110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101111000000;
neuron_parameter[189] <= 368'b11000011100110010001110110101000110110000010101011011000101001111011100010101110111010001100101110101000010111100010100010011010101011000001011110101000100110101010100010000011001010110110101000101011010010101010101010101010101010101010010110110111100111000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101111010000;
neuron_parameter[190] <= 368'b00001010101011111110101010101000001001100000101100010100011010110010010001001010100000001101001110000010110100110000101011010110100010100001001110000100001100111001010100000010000101001010001110111010101010001000000000011001001010101010101001101000111000110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101111100000;
neuron_parameter[191] <= 368'b10001010101101010010101010101000101100001010101101000101000101100001010100101011100110011010101110101001101010100010101010001000001010101001111110101010011011101010101101011111001010100100111110101011010010110011000000101011001000010010100101010011010010000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001101111110000;
neuron_parameter[192] <= 368'b10101010101010000110010110101001110101010001001011010101010101001111000101011010011010100100101100101010000010101010101010101010001010101010101010100010101001101000000000000110100000010111111010011001100010100010000000000011110010101111011011010111000111010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110000000000;
neuron_parameter[193] <= 368'b00101010101010110010000010000100101100100101010110111000000001011001100010101011100100001010100110010000101010011000100001011010101010100100111100101001001010100010100110100100101010101000010010101001010001111010101000010100001010101010110110010010100101100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110000010000;
neuron_parameter[194] <= 368'b01101010101010000110001010101010101100101010101100100010101010110010101010101001101000010101101110010101011100111001010111011010110101000101011010100000010100101010101010000001101010101010101010001010101010101110001010001010101010101010100000011100100001000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110000100000;
neuron_parameter[195] <= 368'b11101010101000111001101000100101100110001010101010111000100010111111001001000001101000101010001010000010101010101000001001001010101000000100001111010100110110101100101011011010101010101101101001010100010010101101010001001010001000101010100100110101110101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110000110000;
neuron_parameter[196] <= 368'b11000010101010001110101010101010101010101010100000100000001010100010100001101010101000000100101110100000011010111011011001101011101000100110101110101010011010111010101100101011001010010010101010101000101010011010010010101001000101011011000001101110000010110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110001000000;
neuron_parameter[197] <= 368'b01110011010100110111010101100101101010101010001000101010101010111010101010101011101010010101101110100101010100101101010010010101101101001001010100010010100100010011010100101000101000010100100100100010100000010011101010101001011010101010110111001101100111010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110001010000;
neuron_parameter[198] <= 368'b01101010101010001010111001111010101100100010101010110010000000111001101001000010101000010101001010001001010100100100010101101010111001010010001101010101000001101001010010010010001101001000101110101100101010111000001011011000101010101010110011011100101100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110001100000;
neuron_parameter[199] <= 368'b01110101011110100101010000010101100101101010101100011000001010100111100010101011101010010010101110101100100000111010110010010111101100010101011110010001010100101010001100101011101000010010101010101001101010101010101010101011001010101010101010011000110010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110001110000;
neuron_parameter[200] <= 368'b10001010101011100110101010101011101010101101001010101010110110110010101011010011100110001101001010001010101100111000101011100010100110100111001010010010011100101001010001110011100011000000101010100100101010111000000010101011001010101010101010100010100111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110010000000;
neuron_parameter[201] <= 368'b10011010101000010110101010011010001000100101001101100011000101101010000100010011101010011010101110101001001010101010101000101010101000100010111110000000011010101011010100100011000101010010101010010100001010101010010010001001101000011010100000010101101100010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110010010000;
neuron_parameter[202] <= 368'b01101010101011101110101010100011010010100101001000001011010100010110100101010101010011010100010100000001000001111110001101101010001010000110101110100001001000101000010100101111001101011010100010110110101110101010001001101011001010101010000000011011101000010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110010100000;
neuron_parameter[203] <= 368'b10001010101010111110101010010111001010100101010010101000000100101010100000100100101010001010010010101100101011001010101000001111101010010010011010110100101011100010011010101000001101001000101110100100000010110010100001000110011010100010100010100100001100000000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110010110000;
neuron_parameter[204] <= 368'b01001010101011110000101010101001001101001010101110110000101000111011001001101001100100010100011011010101001001100001010101010010101001010100111010101000101000101010101010010000111010100101001011001001010100100001000100101000001010111010111101001101110101110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110011000000;
neuron_parameter[205] <= 368'b10001010101010000100011100101100010001110100101101100110010010100001010011001001110000101100001110101110011010101010101100000010101010010110001011101101010010100110110110000011100011011001001001001001110010010101101100101011101010001010101111001000100111100000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001110011010000;
neuron_parameter[206] <= 368'b11101010101001111110101010101000001010101010100100101000101010100100000100100110100110110000101011000010000000111100000110000010010101011001001010010100100000101000001010000111001010101100111110101010010001100010101101000111000010010101010111101010011000010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110011100000;
neuron_parameter[207] <= 368'b10110001101101001010010000000000001010001011001011111010001000100011101001001011100110010101011010010000100101101101011010110100100001001010010010100101000001010010000111100101101010010101010110101011100110010010101010101011101010101010101011110110101010010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110011110000;
neuron_parameter[208] <= 368'b10001010101011010110111100101011000101010010101100011000001010101010010001101010101001010110101111101001001010100110100000100010101010100101011100010000110101101110100011000110001001101111111110100011010010101100100010101010101011101010101110001001101110000000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001110100000000;
neuron_parameter[209] <= 368'b11101111010011111101111000011100100010101011101100001010010010110000101000101010100010111010101010001000101010101010101101001110101011010000101110101101010010101011100101101011100100011010101110100100101010100010101010101010101010101010101010011111101001010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001110100010000;
neuron_parameter[210] <= 368'b11101010101001111010101010101001101010010010110000000001001011111001000001101010100100100110001111011010111101101100101010100111110010101010001000001110100010101011111001000011001010010000001110101001010100100010101000001011101010101010101100011100010010010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110100100000;
neuron_parameter[211] <= 368'b01011010101111000110101000101000111011001010101000101000001010101110001000101010111100100010100110101010001110111011101000101001000110110010111000111011001010101010101100101011101010100010101000101000001010011010111001101010101010010010100100011101101101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110100110000;
neuron_parameter[212] <= 368'b11101010100001110110101010101010001010101010111101001010100001000101000010110011010101011001011001000100010100111100000101000011011000100010101010100010101010101011000010101110101010001010010000100000101001111010000101010001011010100000100100111011111010010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110101000000;
neuron_parameter[213] <= 368'b01101010101010110110000100111000001000001000100010111010010011001001001000001010100100101011100010010100101010011001000010101011001010100100001100101011011011101010100100100110101010001010110010101000010101100010100100010110101010101110100011100111101011100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110101010000;
neuron_parameter[214] <= 368'b01101010101010001000101010000000001010101010101010100010101010111010100010100010100000010101011010101001010101101000100000010111110000010101011110010101010000101001010010100010100100001010001010100010100000100101001010101011101010101010110101001000101100000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110101100000;
neuron_parameter[215] <= 368'b00001010101010100110001010101000101110101000111010101010101110111010100010010011101010000001001010101000010000101010101001000011101010100001001011001000011000101101010101101010110101001010101001001010101010111010101010101001001010101010011101000100110110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110101110000;
neuron_parameter[216] <= 368'b10101010101001111110101010101011101011100010101110100100010010100011010101011010111001000101001011010110100000100000011000000011110001100110001010110010001011111010001010100111101010101101011110010101000101001101010101010101110100010101100101110010011110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110110000000;
neuron_parameter[217] <= 368'b11111100010000010110110101000101001010100011001111101010100010111010100000101010101010000010101100101001000000111011000010101000101010001010100010101000101010010010010101010101101111010101000100101000010101011011101010101000001010101010101110111110111010000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110110010000;
neuron_parameter[218] <= 368'b00101010101010111010101001101010001010100100101111101010100010101010100010001011101000001100101110101000000010101010101100101001101010010010111100100111011010101011001001101011011010100110101011010100101010010100010110101011101011101010111101101100000001100000000000000000000000000011111111110000000011111111111111111010000000000000000000000000000000000001110110100000;
neuron_parameter[219] <= 368'b10100101010110101101010100010101000000110000101000101010000010100110101000101011101000010010101010101100001000100010010010000100101001001001011010100100010101101010010001011011101001100000101010110010010010110010101010101001101010101010011110110010110111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110110110000;
neuron_parameter[220] <= 368'b00001010101011110010101010101001001000010110111010101000011111100000011011010110100000101010011010011010101001110000101010110110110110101010001101001010100010101001001011100011100001000000001110100011000010001010000001101000101010001010100110101000000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110111000000;
neuron_parameter[221] <= 368'b11111010101011111110101110101001101100001000101100010101001100101101010101000011111010010110101110101011000010100010101000101011101010110011011010101101011010101011110000001010000110001011011110010000001000011001000100011000101000100010101011100110101100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001110111010000;
neuron_parameter[222] <= 368'b10101010101010010010101110100000110010110101001111001001110011101100100100110101010011010110000101001101011011111100000101101011011010000110101010110010101010101010100101101010101000010100111010100101001000111010010100100001101000011000110100111011110011010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001110111100000;
neuron_parameter[223] <= 368'b10101010101010011010100001010110101010010101010110100000101101001010010010101100101010001010110110101001010010001010101101001011101010100010101010110010101011001011010010010000101010110101011110100000010011101010101010101100101010101010101100001000000110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001110111110000;
neuron_parameter[224] <= 368'b10001010101011101110101010101010010011100001001100001110101010111010101000101010101010100010101010101001000000110001010100010110101100111101001110100000110110101011001011101010100110100110011010011010111101101001111010011001101010101010101001011110111001100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111000000000;
neuron_parameter[225] <= 368'b11001010101001010001011100101101010101010000111101000001101000111101010101100001100000001010111010100000101011110010001001100010111010110101011011001011010000111100100100001010110010110100001001001010010100111100001011000001101011101010101101100000100101000000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001111000010000;
neuron_parameter[226] <= 368'b10001010101100010110101010101011101000111010101110100001010110100011010101010011110001001000001110000001101000111001100100101010100010010100001110000000000001101010101010000111101010101001011111010101000101110001010101010101010101010101000000010110001000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111000100000;
neuron_parameter[227] <= 368'b01111001001101111111100010101101101010101001011110101000010101100010100101001111101101011010111010010100101101110000010010100001101011011010110010111001011011010010010101100100101000010010000110100000101000011010101010101010101010101010100110110000111100000000000000000000000000000011111111110000000011111111110000000100000000000000000000000000000000000001111000110000;
neuron_parameter[228] <= 368'b11101010101010100110110101101011000111010100101100101001001000100000000010101010100000001010101110000101010000100010010101011011111010110100001001001010010101101010001001010110001010100100001110110000010110110100101010011001101010101010100110000110100110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111001000000;
neuron_parameter[229] <= 368'b00100101010110010001010101010110000101001011101110100100000010110010100010100010111001101010101000101000101010110010000010101110101001001001011110100100110101101011110101010110101001010010101010101000000010110010101010101001101010101010111010100100110000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111001010000;
neuron_parameter[230] <= 368'b00001010101010010110101010101011101010110110001110101010110100111010000010001011101001101011001110010010100100111001001010000010100110101001101000010010100000101001001010100011000101101010001110110100000010100010100110101000101010101010100100101010001111100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111001100000;
neuron_parameter[231] <= 368'b11001010101011100110101010111010011001000101001000100100100101101110100010101011111010110000101010101011001010110000100101001010000011010001011010011001001011101010000100101011001100001010111110000010101010101011101010011001001010101010100100010001100000110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111001110000;
neuron_parameter[232] <= 368'b11001010101011011010101010101011000101101010001011010100100101001011000010010010011010101101001001101000010100110101001001000010010000100010101010010010101010101000001010101010111001000010100110110100101010110110010101010000011010100101001111001111111011110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111010000000;
neuron_parameter[233] <= 368'b00101010101010000010001101010110001010001011010010101000001000111010110010010100101001000010010010100010000001000010100000100010001001011010101110100100101001001001011010010111101101100101101010010110100010111010010010110111101010000010100101011100100000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111010010000;
neuron_parameter[234] <= 368'b11101010101010101110100010110010001010001000101010101010101010101010100000010110101000010001011010100100100101100001000001010111101100010101011111110001010010101001000010101010100100101010001010100010101010110000000010101000001010101010101111001100101010000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001111010100000;
neuron_parameter[235] <= 368'b00101010101000110001010101001100101101010110001110010000000001111000010010101001110100101010101000011010000010111000001000001011101000101101001010101010110000100110101011010010110100000100101101010100110000101101100011011001101100101010111100011100100110100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001111010110000;
neuron_parameter[236] <= 368'b01001010101010100110101010101011101001101010100100110011000010110011000101001011110110100000101011001011010110110101001101011011110110110101101010101011110010101010101100101010101010110010101111000010101010010101000001000010110101010101010010011100001110000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111011000000;
neuron_parameter[237] <= 368'b01010101010001000011101101000101001010101101001100100010110000110010001011101011101100100110101100101010101000110000001010100001100000101001010100100100110101010011010010101001000100010100100110101010011000010010101010101000011010101010100010101100011010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111011010000;
neuron_parameter[238] <= 368'b00001010101010011110100110101011100011010010101000111000001010101011100000011010101000110100101011101001011000101010100101101011100000110101101001010001010111101101001101010111010010100010111010001011001010111010101111101001001010101010111101101000100100110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111011100000;
neuron_parameter[239] <= 368'b01000110111010101111101010101001100000101011001000001000111010101000100011101011100010000101001010000100010111111001010101000010100100010110011010110001001001101010100100100011111010010010101010101001010010100010101100101000001010101010101101000001101110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111011110000;
neuron_parameter[240] <= 368'b01101010101010010010101010101011001010000101111100101000010100111001000001010110100000001000011011010010101000100101001010001011110101000100001010000101010001101010100010010011001010111100101110011101010000110000110101101000001010101010100101001000100001100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001111100000000;
neuron_parameter[241] <= 368'b10001010101011110010101110101011011001010010001001010101100001110101010000101010111100100110101110101011010010111010101000001011101010011011011010110100110011101011110100001111101011010101111110101000010100100000001010001000001000110010001101100101110110110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001111100010000;
neuron_parameter[242] <= 368'b10101010101011011110111010101000111100101001001001010110110001000100001011010110010100110100101001001001010010111110101010101011011011101010101110111100100000111000110101000110101110110110010010110010010010100010011010000000011010101000000110001011111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111100100000;
neuron_parameter[243] <= 368'b01001010101000100110001101111010001110001000110000111000000011100001010000000011100100101010100010010110101010000001000010000010101010100100001100101011011011100010100100100111001010001010011010101000110101111010101000010100011010101010100111001101101100010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001111100110000;
neuron_parameter[244] <= 368'b11101010101011000000101010101000101110101010101100110000001010110011100100101000100101101110101010010100110110101101010001011111111100010101111010100101010001001010000000010010110010101001001010001010101010011111001000101011101010101010111000101010100110010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001111101000000;
neuron_parameter[245] <= 368'b10101010101010011001010101101011110110101111111100001100001110101010110000001011101010011010001110101010000000111010100101010010101010110110101011001010011010100101010001101011110100001110101101001010111010101010101011101000001000101010110101100110100000110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001111101010000;
neuron_parameter[246] <= 368'b10001010101001001010101010101000001000000010100110110001010010111111001011011011100000101101101010111010110110101011101011011010100110101101101110101010010010101010100101101011101010000010101010110100101010011001010110101010010101011111011011010110001100100000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001111101100000;
neuron_parameter[247] <= 368'b00111000101000100111101000010100001010000101011000101000001101111010000000101010100101101010111110110100101010100000010110101001101010010100100110110101000100010011010001010001100010010101100110101001010010010010101010101011101010101010100101101000110101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001111101110000;
neuron_parameter[248] <= 368'b00001010101011000010010110101011001110010010101110101000011010100010110001001010101010010110101110101001001010110000101000101010100100101101001001011010100111101110111010110111001110110111001110000011101010100100011010101000101010101010101101111001101110010000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001111110000000;
neuron_parameter[249] <= 368'b11100001011010000101100001011110000110101011101000011010000010110101101000101010101010111010101000111001101011100010100001101110101010010110101010111000011010101011000001101010101100001010101010101100101010000010101010101000001010101010100010101101110010110000000000000000000000000011111111110000000011111111111111111100000000000000000000000000000000000001111110010000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                neuron_parameter[neuron_num][111:103] <= potential_out;
            end
        end
    end
    else begin
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
                neuron_parameter[0] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[1] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[2] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[3] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[4] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[5] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[6] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[7] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[8] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[9] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[10] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[11] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[12] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[13] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[14] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[15] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[16] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[17] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[18] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[19] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[20] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[21] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[22] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[23] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[24] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[25] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[26] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[27] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[28] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[29] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[30] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[31] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[32] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[33] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[34] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[35] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[36] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[37] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[38] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[39] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[40] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[41] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[42] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[43] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[44] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[45] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[46] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[47] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[48] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[49] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[50] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[51] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[52] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[53] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[54] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[55] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[56] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[57] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[58] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[59] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[60] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[61] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[62] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[63] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
            end
            else if(update_potential) begin
                neuron_parameter[neuron_num][111:103] <= potential_out;
            end
        end
    end
endgenerate

assign neuron_instructions[0] = 2'b00;
assign neuron_instructions[1] = 2'b01;
assign neuron_instructions[2] = 2'b00;
assign neuron_instructions[3] = 2'b01;
assign neuron_instructions[4] = 2'b00;
assign neuron_instructions[5] = 2'b01;
assign neuron_instructions[6] = 2'b00;
assign neuron_instructions[7] = 2'b01;
assign neuron_instructions[8] = 2'b00;
assign neuron_instructions[9] = 2'b01;
assign neuron_instructions[10] = 2'b00;
assign neuron_instructions[11] = 2'b01;
assign neuron_instructions[12] = 2'b00;
assign neuron_instructions[13] = 2'b01;
assign neuron_instructions[14] = 2'b00;
assign neuron_instructions[15] = 2'b01;
assign neuron_instructions[16] = 2'b00;
assign neuron_instructions[17] = 2'b01;
assign neuron_instructions[18] = 2'b00;
assign neuron_instructions[19] = 2'b01;
assign neuron_instructions[20] = 2'b00;
assign neuron_instructions[21] = 2'b01;
assign neuron_instructions[22] = 2'b00;
assign neuron_instructions[23] = 2'b01;
assign neuron_instructions[24] = 2'b00;
assign neuron_instructions[25] = 2'b01;
assign neuron_instructions[26] = 2'b00;
assign neuron_instructions[27] = 2'b01;
assign neuron_instructions[28] = 2'b00;
assign neuron_instructions[29] = 2'b01;
assign neuron_instructions[30] = 2'b00;
assign neuron_instructions[31] = 2'b01;
assign neuron_instructions[32] = 2'b00;
assign neuron_instructions[33] = 2'b01;
assign neuron_instructions[34] = 2'b00;
assign neuron_instructions[35] = 2'b01;
assign neuron_instructions[36] = 2'b00;
assign neuron_instructions[37] = 2'b01;
assign neuron_instructions[38] = 2'b00;
assign neuron_instructions[39] = 2'b01;
assign neuron_instructions[40] = 2'b00;
assign neuron_instructions[41] = 2'b01;
assign neuron_instructions[42] = 2'b00;
assign neuron_instructions[43] = 2'b01;
assign neuron_instructions[44] = 2'b00;
assign neuron_instructions[45] = 2'b01;
assign neuron_instructions[46] = 2'b00;
assign neuron_instructions[47] = 2'b01;
assign neuron_instructions[48] = 2'b00;
assign neuron_instructions[49] = 2'b01;
assign neuron_instructions[50] = 2'b00;
assign neuron_instructions[51] = 2'b01;
assign neuron_instructions[52] = 2'b00;
assign neuron_instructions[53] = 2'b01;
assign neuron_instructions[54] = 2'b00;
assign neuron_instructions[55] = 2'b01;
assign neuron_instructions[56] = 2'b00;
assign neuron_instructions[57] = 2'b01;
assign neuron_instructions[58] = 2'b00;
assign neuron_instructions[59] = 2'b01;
assign neuron_instructions[60] = 2'b00;
assign neuron_instructions[61] = 2'b01;
assign neuron_instructions[62] = 2'b00;
assign neuron_instructions[63] = 2'b01;
assign neuron_instructions[64] = 2'b00;
assign neuron_instructions[65] = 2'b01;
assign neuron_instructions[66] = 2'b00;
assign neuron_instructions[67] = 2'b01;
assign neuron_instructions[68] = 2'b00;
assign neuron_instructions[69] = 2'b01;
assign neuron_instructions[70] = 2'b00;
assign neuron_instructions[71] = 2'b01;
assign neuron_instructions[72] = 2'b00;
assign neuron_instructions[73] = 2'b01;
assign neuron_instructions[74] = 2'b00;
assign neuron_instructions[75] = 2'b01;
assign neuron_instructions[76] = 2'b00;
assign neuron_instructions[77] = 2'b01;
assign neuron_instructions[78] = 2'b00;
assign neuron_instructions[79] = 2'b01;
assign neuron_instructions[80] = 2'b00;
assign neuron_instructions[81] = 2'b01;
assign neuron_instructions[82] = 2'b00;
assign neuron_instructions[83] = 2'b01;
assign neuron_instructions[84] = 2'b00;
assign neuron_instructions[85] = 2'b01;
assign neuron_instructions[86] = 2'b00;
assign neuron_instructions[87] = 2'b01;
assign neuron_instructions[88] = 2'b00;
assign neuron_instructions[89] = 2'b01;
assign neuron_instructions[90] = 2'b00;
assign neuron_instructions[91] = 2'b01;
assign neuron_instructions[92] = 2'b00;
assign neuron_instructions[93] = 2'b01;
assign neuron_instructions[94] = 2'b00;
assign neuron_instructions[95] = 2'b01;
assign neuron_instructions[96] = 2'b00;
assign neuron_instructions[97] = 2'b01;
assign neuron_instructions[98] = 2'b00;
assign neuron_instructions[99] = 2'b01;
assign neuron_instructions[100] = 2'b00;
assign neuron_instructions[101] = 2'b01;
assign neuron_instructions[102] = 2'b00;
assign neuron_instructions[103] = 2'b01;
assign neuron_instructions[104] = 2'b00;
assign neuron_instructions[105] = 2'b01;
assign neuron_instructions[106] = 2'b00;
assign neuron_instructions[107] = 2'b01;
assign neuron_instructions[108] = 2'b00;
assign neuron_instructions[109] = 2'b01;
assign neuron_instructions[110] = 2'b00;
assign neuron_instructions[111] = 2'b01;
assign neuron_instructions[112] = 2'b00;
assign neuron_instructions[113] = 2'b01;
assign neuron_instructions[114] = 2'b00;
assign neuron_instructions[115] = 2'b01;
assign neuron_instructions[116] = 2'b00;
assign neuron_instructions[117] = 2'b01;
assign neuron_instructions[118] = 2'b00;
assign neuron_instructions[119] = 2'b01;
assign neuron_instructions[120] = 2'b00;
assign neuron_instructions[121] = 2'b01;
assign neuron_instructions[122] = 2'b00;
assign neuron_instructions[123] = 2'b01;
assign neuron_instructions[124] = 2'b00;
assign neuron_instructions[125] = 2'b01;
assign neuron_instructions[126] = 2'b00;
assign neuron_instructions[127] = 2'b01;
assign neuron_instructions[128] = 2'b00;
assign neuron_instructions[129] = 2'b01;
assign neuron_instructions[130] = 2'b00;
assign neuron_instructions[131] = 2'b01;
assign neuron_instructions[132] = 2'b00;
assign neuron_instructions[133] = 2'b01;
assign neuron_instructions[134] = 2'b00;
assign neuron_instructions[135] = 2'b01;
assign neuron_instructions[136] = 2'b00;
assign neuron_instructions[137] = 2'b01;
assign neuron_instructions[138] = 2'b00;
assign neuron_instructions[139] = 2'b01;
assign neuron_instructions[140] = 2'b00;
assign neuron_instructions[141] = 2'b01;
assign neuron_instructions[142] = 2'b00;
assign neuron_instructions[143] = 2'b01;
assign neuron_instructions[144] = 2'b00;
assign neuron_instructions[145] = 2'b01;
assign neuron_instructions[146] = 2'b00;
assign neuron_instructions[147] = 2'b01;
assign neuron_instructions[148] = 2'b00;
assign neuron_instructions[149] = 2'b01;
assign neuron_instructions[150] = 2'b00;
assign neuron_instructions[151] = 2'b01;
assign neuron_instructions[152] = 2'b00;
assign neuron_instructions[153] = 2'b01;
assign neuron_instructions[154] = 2'b00;
assign neuron_instructions[155] = 2'b01;
assign neuron_instructions[156] = 2'b00;
assign neuron_instructions[157] = 2'b01;
assign neuron_instructions[158] = 2'b00;
assign neuron_instructions[159] = 2'b01;
assign neuron_instructions[160] = 2'b00;
assign neuron_instructions[161] = 2'b01;
assign neuron_instructions[162] = 2'b00;
assign neuron_instructions[163] = 2'b01;
assign neuron_instructions[164] = 2'b00;
assign neuron_instructions[165] = 2'b01;
assign neuron_instructions[166] = 2'b00;
assign neuron_instructions[167] = 2'b01;
assign neuron_instructions[168] = 2'b00;
assign neuron_instructions[169] = 2'b01;
assign neuron_instructions[170] = 2'b00;
assign neuron_instructions[171] = 2'b01;
assign neuron_instructions[172] = 2'b00;
assign neuron_instructions[173] = 2'b01;
assign neuron_instructions[174] = 2'b00;
assign neuron_instructions[175] = 2'b01;
assign neuron_instructions[176] = 2'b00;
assign neuron_instructions[177] = 2'b01;
assign neuron_instructions[178] = 2'b00;
assign neuron_instructions[179] = 2'b01;
assign neuron_instructions[180] = 2'b00;
assign neuron_instructions[181] = 2'b01;
assign neuron_instructions[182] = 2'b00;
assign neuron_instructions[183] = 2'b01;
assign neuron_instructions[184] = 2'b00;
assign neuron_instructions[185] = 2'b01;
assign neuron_instructions[186] = 2'b00;
assign neuron_instructions[187] = 2'b01;
assign neuron_instructions[188] = 2'b00;
assign neuron_instructions[189] = 2'b01;
assign neuron_instructions[190] = 2'b00;
assign neuron_instructions[191] = 2'b01;
assign neuron_instructions[192] = 2'b00;
assign neuron_instructions[193] = 2'b01;
assign neuron_instructions[194] = 2'b00;
assign neuron_instructions[195] = 2'b01;
assign neuron_instructions[196] = 2'b00;
assign neuron_instructions[197] = 2'b01;
assign neuron_instructions[198] = 2'b00;
assign neuron_instructions[199] = 2'b01;
assign neuron_instructions[200] = 2'b00;
assign neuron_instructions[201] = 2'b01;
assign neuron_instructions[202] = 2'b00;
assign neuron_instructions[203] = 2'b01;
assign neuron_instructions[204] = 2'b00;
assign neuron_instructions[205] = 2'b01;
assign neuron_instructions[206] = 2'b00;
assign neuron_instructions[207] = 2'b01;
assign neuron_instructions[208] = 2'b00;
assign neuron_instructions[209] = 2'b01;
assign neuron_instructions[210] = 2'b00;
assign neuron_instructions[211] = 2'b01;
assign neuron_instructions[212] = 2'b00;
assign neuron_instructions[213] = 2'b01;
assign neuron_instructions[214] = 2'b00;
assign neuron_instructions[215] = 2'b01;
assign neuron_instructions[216] = 2'b00;
assign neuron_instructions[217] = 2'b01;
assign neuron_instructions[218] = 2'b00;
assign neuron_instructions[219] = 2'b01;
assign neuron_instructions[220] = 2'b00;
assign neuron_instructions[221] = 2'b01;
assign neuron_instructions[222] = 2'b00;
assign neuron_instructions[223] = 2'b01;
assign neuron_instructions[224] = 2'b00;
assign neuron_instructions[225] = 2'b01;
assign neuron_instructions[226] = 2'b00;
assign neuron_instructions[227] = 2'b01;
assign neuron_instructions[228] = 2'b00;
assign neuron_instructions[229] = 2'b01;
assign neuron_instructions[230] = 2'b00;
assign neuron_instructions[231] = 2'b01;
assign neuron_instructions[232] = 2'b00;
assign neuron_instructions[233] = 2'b01;
assign neuron_instructions[234] = 2'b00;
assign neuron_instructions[235] = 2'b01;
assign neuron_instructions[236] = 2'b00;
assign neuron_instructions[237] = 2'b01;
assign neuron_instructions[238] = 2'b00;
assign neuron_instructions[239] = 2'b01;
assign neuron_instructions[240] = 2'b00;
assign neuron_instructions[241] = 2'b01;
assign neuron_instructions[242] = 2'b00;
assign neuron_instructions[243] = 2'b01;
assign neuron_instructions[244] = 2'b00;
assign neuron_instructions[245] = 2'b01;
assign neuron_instructions[246] = 2'b00;
assign neuron_instructions[247] = 2'b01;
assign neuron_instructions[248] = 2'b00;
assign neuron_instructions[249] = 2'b01;
assign neuron_instructions[250] = 2'b00;
assign neuron_instructions[251] = 2'b01;
assign neuron_instructions[252] = 2'b00;
assign neuron_instructions[253] = 2'b01;
assign neuron_instructions[254] = 2'b00;
assign neuron_instructions[255] = 2'b01;

endmodule
